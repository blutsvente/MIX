        /* ------------------------------------------------------------
          Generator information:
          used package Micronas::Reg is version 1.88  
          this package RegViews.pm is version 1.93
          use with RTL libraries (this release or higher):
          ip_ocp/0002/ip_ocp_016_21Jan2009
          ip_sync/0001/ip_sync_006_23jan2008
        ------------------------------------------------------------ */

// useful defines for domain fe1
`define cvbsdetect_msb_c  'h02
`define dgatel_msb_c      'h03
`define dgates_msb_c      'h04
`define dummy_fe_msb_c    'h02
`define mvstart_msb_c     'h03
`define mvstop_msb_c      'h03
`define r_test_msb_c      'h02
`define reg_0x0_offs_c    'h0000
`define reg_0x10_offs_c   'h0010
`define reg_0x14_offs_c   'h0014
`define reg_0x18_offs_c   'h0018
`define reg_0x1C_offs_c   'h001c
`define reg_0x20_offs_c   'h0020
`define reg_0x28_offs_c   'h0028
`define reg_0x4_offs_c    'h0004
`define reg_0x8_offs_c    'h0008
`define reg_0xC_offs_c    'h000c
`define sha_r_test_msb_c  'h07
`define sha_rw2_msb_c     'h1f
`define sha_w_test_msb_c  'h03
`define usr_ali_msb_c     'h01
`define usr_rw_test_msb_c 'h03
`define usr_w_test_msb_c  'h03
`define w_test_msb_c      'h03
`define wd_16_test2_msb_c 'h07
`define wd_16_test_msb_c  'h0f
// end
