-- -------------------------------------------------------------
--
-- Generated Architecture Declaration for rtl of ent_b
--
-- Generated
--  by:  wig
--  on:  Thu Jun 29 16:41:09 2006
--  cmd: /cygdrive/h/work/eclipse/MIX/mix_0.pl -conf macro._MP_VHDL_USE_ENTY_MP_=Overwritten vhdl_enty from cmdline -conf macro._MP_VHDL_HOOK_ARCH_BODY_MP_=Use macro vhdl_hook_arch_body -conf macro._MP_ADD_MY_OWN_MP_=overloading my own macro ../../configuration.xls
--
-- !!! Do not edit this file! Autogenerated by MIX !!!
-- $Author: wig $
-- $Id: ent_b-rtl-a.vhd,v 1.1 2006/07/04 09:54:10 wig Exp $
-- $Date: 2006/07/04 09:54:10 $
-- $Log: ent_b-rtl-a.vhd,v $
-- Revision 1.1  2006/07/04 09:54:10  wig
-- Update more testcases, add configuration/cfgfile
--
--
-- Based on Mix Architecture Template built into RCSfile: MixWriter.pm,v 
-- Id: MixWriter.pm,v 1.90 2006/06/22 07:13:21 wig Exp 
--
-- Generator: mix_0.pl Revision: 1.46 , wilfried.gaensheimer@micronas.com
-- (C) 2003,2005 Micronas GmbH
--
-- --------------------------------------------------------------
-- modifiy vhdl_use_arch 
library IEEE;
use IEEE.std_logic_1164.all;

-- No project specific VHDL libraries/arch

typedef vhdl_use_arch_def std_ulogic_vector;
-- end of vhdl_use_arch

--
--
-- Start of Generated Architecture rtl of ent_b
--
architecture rtl of ent_b is 

	--
	-- Generated Constant Declarations
	--


	--
	-- Generated Components
	--
	component ent_ba
		-- No Generated Generics
		-- No Generated Port
	end component;
	-- ---------

	component ent_bb
		-- No Generated Generics
		-- No Generated Port
	end component;
	-- ---------



	--
	-- Generated Signal List
	--
	--
	-- End of Generated Signal List
	--




begin

Use macro vhdl_hook_arch_body
	--
	-- Generated Concurrent Statements
	--

	--
	-- Generated Signal Assignments
	--


	--
	-- Generated Instances and Port Mappings
	--
		-- Generated Instance Port Map for inst_ba
		inst_ba: ent_ba

		;

		-- End of Generated Instance Port Map for inst_ba

		-- Generated Instance Port Map for inst_bb
		inst_bb: ent_bb

		;

		-- End of Generated Instance Port Map for inst_bb



end rtl;


--
--!End of Architecture/s
-- --------------------------------------------------------------
