 a @          :           Telex/     Telex   b @          ,:           ISDN0     ISDN   c @          -:           TTYTDD1     TTYTDD   d @          K:           
OtherPhone2     
OtherPhone   l @          :           OtherFax3     OtherFax   n @          #:           CompanyMainPhone4     CompanyMainPhone   ` @          W:           PrimaryPhone5     PrimaryPhone   | @          :           CallbackPhone6     CallbackPhone   { @          :           Private7     Private     @          6           
Profession;   "  
Profession   Y @          F:           NickName8     NickName   \ @          O:           ManagerName9      ManagerName   X @          N:           
ReferredBy:   !  
ReferredBy   y @          G:           Hobbies<   #  Hobbies   r @          C:           Account=   $  Account   x @           :           FTPSite>   %  FTPSite   s @          L:           PersonalHomePage?   &  PersonalHomePage   U @          P:           Mileage@   '  Mileage   �  @&{00062008-0000-0000-C000-000000000046} 4�      F�           BillingInformationA   (  BillingInformation   �  @&{00062008-0000-0000-C000-000000000046} 5�      G�           OrganizationalIdNumberB   )  OrganizationalIdNumber   �  @          