        /* ------------------------------------------------------------
          Generator information:
          used package Micronas::Reg is version 1.90  
          package RegViewURAC is version 1.3
          use with RTL libraries (this release or higher):
          ip_sync/0001/ip_sync_006_23jan2008
        ------------------------------------------------------------ */

// useful defines for domain urac_fe1
`define FE_MVDET_offs_c       'h03
`define FE_NATIVE_offs_c      'h04
`define FE_NT_offs_c          'h05
`define FE_YCDET_CTRL2_offs_c 'h02
`define FE_YCDET_CTRL_offs_c  'h00
`define FE_YCDET_STAT_offs_c  'h01
`define cvbsdetect2_pos_c     'h0
`define cvbsdetect2_size_c    'h1
`define cvbsdetect_pos_c      'h0
`define cvbsdetect_size_c     'h1
`define dgatel_lsb_c          'h0
`define dgatel_msb_c          'h3
`define dgatel_pos_c          'h0
`define dgatel_size_c         'h4
`define dgates_lsb_c          'h0
`define dgates_msb_c          'h3
`define dgates_pos_c          'h4
`define dgates_size_c         'h4
`define mvstart_lsb_c         'h0
`define mvstart_msb_c         'h4
`define mvstart_pos_c         'h0
`define mvstart_size_c        'h5
`define mvstop_lsb_c          'h0
`define mvstop_msb_c          'h2
`define mvstop_pos_c          'h5
`define mvstop_size_c         'h3
`define prova_lsb_c           'h0
`define prova_msb_c           'h4
`define prova_pos_c           'h0
`define prova_size_c          'h5
`define r_native_lsb_c        'h0
`define r_native_msb_c        'h1
`define r_native_pos_c        'h2
`define r_native_size_c       'h2
`define rw_native_lsb_c       'h0
`define rw_native_msb_c       'h1
`define rw_native_pos_c       'h0
`define rw_native_size_c      'h2
`define y_test_pos_c          'h2
`define y_test_size_c         'h1
`define ycdetect2_pos_c       'h1
`define ycdetect2_size_c      'h1
`define ycdetect_pos_c        'h1
`define ycdetect_size_c       'h1
// end
