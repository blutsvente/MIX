        /* ------------------------------------------------------------
          Generator information:
          used package Micronas::Reg is version 1.96  
          package RegViewIHB is version 1.6
          use with RTL libraries (this release or higher):
          ip_ocp/0002/ip_ocp_018_13Feb2009
          ip_sync/0001/ip_sync_006_23jan2008
        ------------------------------------------------------------ */

// useful defines for domain fe1
`define cvbsdetect_lsb_c   'h00
`define cvbsdetect_msb_c   'h02
`define cvbsdetect_pos_c   'h00
`define cvbsdetect_size_c  'h03
`define dgatel_lsb_c       'h00
`define dgatel_msb_c       'h03
`define dgatel_pos_c       'h00
`define dgatel_size_c      'h04
`define dgates_lsb_c       'h00
`define dgates_msb_c       'h04
`define dgates_pos_c       'h04
`define dgates_size_c      'h05
`define dummy_fe_lsb_c     'h00
`define dummy_fe_msb_c     'h02
`define dummy_fe_pos_c     'h09
`define dummy_fe_size_c    'h03
`define mvstart_lsb_c      'h00
`define mvstart_msb_c      'h03
`define mvstart_pos_c      'h00
`define mvstart_size_c     'h04
`define mvstop_lsb_c       'h00
`define mvstop_msb_c       'h03
`define mvstop_pos_c       'h04
`define mvstop_size_c      'h04
`define r_test_lsb_c       'h00
`define r_test_msb_c       'h02
`define r_test_pos_c       'h00
`define r_test_size_c      'h03
`define reg_0x0_offs_c     'h0000
`define reg_0x10_offs_c    'h0010
`define reg_0x14_offs_c    'h0014
`define reg_0x18_offs_c    'h0018
`define reg_0x1C_offs_c    'h001c
`define reg_0x20_offs_c    'h0020
`define reg_0x28_offs_c    'h0028
`define reg_0x4_offs_c     'h0004
`define reg_0x8_offs_c     'h0008
`define reg_0xC_offs_c     'h000c
`define sha_r_test_lsb_c   'h00
`define sha_r_test_msb_c   'h07
`define sha_r_test_pos_c   'h03
`define sha_r_test_size_c  'h08
`define sha_rw2_lsb_c      'h00
`define sha_rw2_msb_c      'h1f
`define sha_rw2_pos_c      'h00
`define sha_rw2_size_c     'h20
`define sha_w_test_lsb_c   'h00
`define sha_w_test_msb_c   'h03
`define sha_w_test_pos_c   'h14
`define sha_w_test_size_c  'h04
`define usr_ali_lsb_c      'h00
`define usr_ali_msb_c      'h01
`define usr_ali_pos_c      'h08
`define usr_ali_size_c     'h02
`define usr_r_test_pos_c   'h02
`define usr_r_test_size_c  'h01
`define usr_rw_test_lsb_c  'h00
`define usr_rw_test_msb_c  'h03
`define usr_rw_test_pos_c  'h0b
`define usr_rw_test_size_c 'h04
`define usr_w_test_lsb_c   'h00
`define usr_w_test_msb_c   'h03
`define usr_w_test_pos_c   'h00
`define usr_w_test_size_c  'h04
`define w_test_lsb_c       'h00
`define w_test_msb_c       'h03
`define w_test_pos_c       'h10
`define w_test_size_c      'h04
`define wd_16_test2_lsb_c  'h00
`define wd_16_test2_msb_c  'h07
`define wd_16_test2_pos_c  'h00
`define wd_16_test2_size_c 'h08
`define wd_16_test_lsb_c   'h00
`define wd_16_test_msb_c   'h0f
`define wd_16_test_pos_c   'h00
`define wd_16_test_size_c  'h10
`define ycdetect_pos_c     'h01
`define ycdetect_size_c    'h01
// end
