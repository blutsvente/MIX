-- -------------------------------------------------------------
--
--  Entity Declaration for ent_a
--
-- Generated
--  by:  wig
--  on:  Thu Mar 16 07:48:49 2006
--  cmd: /cygdrive/h/work/eclipse/MIX/mix_0.pl -conf macro._MP_VHDL_USE_ENTY_MP_=Overwritten vhdl_enty from cmdline -conf macro._MP_VHDL_HOOK_ARCH_BODY_MP_=Use macro vhdl_hook_arch_body -conf macro._MP_ADD_MY_OWN_MP_=overloading my own macro -nodelta ../../configuration.xls
--
-- !!! Do not edit this file! Autogenerated by MIX !!!
-- $Author: wig $
-- $Id: ent_a-e.vhd,v 1.1 2006/03/16 14:12:14 wig Exp $
-- $Date: 2006/03/16 14:12:14 $
-- $Log: ent_a-e.vhd,v $
-- Revision 1.1  2006/03/16 14:12:14  wig
-- Added testcase for command line -conf add/overload
--
--
-- Based on Mix Entity Template built into RCSfile: MixWriter.pm,v 
-- Id: MixWriter.pm,v 1.77 2006/03/14 08:10:34 wig Exp 
--
-- Generator: mix_0.pl Version: Revision: 1.44 , wilfried.gaensheimer@micronas.com
-- (C) 2003,2005 Micronas GmbH
--
-- --------------------------------------------------------------
-- adding to vhdl_use_enty
library IEEE;
use IEEE.std_logic_1164.all;

-- Generated use statements
library wig;
use wig.test.all;

typedef use_enty_private std_ulogic_vector;

--

--
-- Start of Generated Entity ent_a
--
entity ent_a is

	-- Generics:
		-- No Generated Generics for Entity ent_a

	-- Generated Port Declaration:
		port(
		-- Generated Port for Entity ent_a
			p_mix_sig_01_go	: out	std_ulogic;
			p_mix_sig_03_go	: out	std_ulogic;
			p_mix_sig_04_gi	: in	std_ulogic;
			p_mix_sig_05_2_1_go	: out	std_ulogic_vector(1 downto 0);
			p_mix_sig_06_gi	: in	std_ulogic_vector(3 downto 0);
			p_mix_sig_i_ae_gi	: in	std_ulogic_vector(6 downto 0);
			p_mix_sig_o_ae_go	: out	std_ulogic_vector(7 downto 0);
			port_i_a	: in	std_ulogic;	-- Input Port
			port_o_a	: out	std_ulogic;	-- Output Port
			sig_07	: in	std_ulogic_vector(5 downto 0);	-- Conflicting definition, IN false!
			sig_08	: out	std_ulogic_vector(8 downto 2);	-- VHDL intermediate needed (port name)
			sig_13	: out	std_ulogic_vector(4 downto 0);	-- Create internal signal name
			sig_i_a2	: in	std_ulogic;	-- Input Port
			sig_o_a2	: out	std_ulogic	-- Output Port
		-- End of Generated Port for Entity ent_a
		);
end ent_a;
--
-- End of Generated Entity ent_a
--


--
--!End of Entity/ies
-- --------------------------------------------------------------
