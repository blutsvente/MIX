��p�e��g��CU��Aq�i�F�6�F��z�u��{�6Q�Q�G�b��Y�!pŘH&l���GQ6h#���.�9k
E�a�� X���J�� �}	}U�QQ��Ѐg<��,��3�rzy�G
�&��/���\���\�������`sD/�HY�9/;<�g�Evn��L�V�����K,�U�:J[���y�-���^p^��C?�zȥ�t�0Ѽ�H}!��mPN�艜Nm���"�3����I�ޛ;�:��8�}+�pAaV��,L*�P�D]��6,GA�AH_6�rOq��� 5n��,EH��x�#�i���*d�ǳ��$!}�Q7����X�}GK�+Ì�M�ߺ˛��W̮�5��1�ūc'���g<�!(�;��6AA$bAA�6A66HA�b�b������E�.��sS �Ε�Я��+�2zz� ̂��-��SA����w�+�Bˢ���j&{63�"���5��&�2��C�՝�M���Qbe��3��e��;�(�O��{+
8ڤ<���b���΃B�A����;~��c4d�+̥1O���8z��E�U{�"����#�A9c�)��k�fx�ӫ��,sD%{*�E)uw3�^�3@d�~�-9�<�-����+'�X&���&�JXP�k%c���e��W=z�J6��•�ZФ�O�]eqi'���t��튕� �3X �B����j
^(yF�1@*����	dc��NTe#-�a�60�����˹��G�հ[Ve?���w�hߠ
�Qg��L=I�����~Ŭk(�7Mz�%u�d��/:�_Y}�����!m����������??�<_�>�:�G{q�H�8��|�~qh g�"�ڪ���j
�BtJ���̲=,�F/D��H&�==========AAAAbAA�6A66HA	A�S========�0=��*�b�����C3|�Y:"�S@���Cn7 A�柰eY�.YS��>�d��E�H�*�0����'AAf6�	6A�A'	AAAbAA�6A66HAYb�n Ak�*n����A���@�A�Х��^�@�v9���w�5+k,`�� �M�Zw���붎;��~��${�G��a��!C��g�6j.S��[��ʷ�4������!��&S����E+�&�"����/�@^�F�<�=���H�q)�Ύ�(Z���C�Re�1�X�[b�]�K3sH0���en]Ƶ��+���$��R��A��γ3NDbg�u�X<���0�1��.�@e�,�]��O�[�����9v���{��v\n��"����Xk��ʾ�����S*n�c�����6�y?����